`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/03/23 00:11:45
// Design Name: 
// Module Name: flush_ctrl
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include	"D:\Grade2\RISC_V\CPU\CPU.srcs\sources_1\config.v"
module flush_ctrl(

    );
endmodule

`timescale 1ns / 1ps
module uart_tb(
    );

reg clk;
reg rst;
reg rx;

wire flag;
wire[31:0] data;
wire[15:0] addr;

initial begin
    clk = 0;
    rst = 1;
    rx = 1;
    #1 
    rst = 0;
    #20.5
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;

    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;

        #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;


    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;


    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;
    #5208
    #5208
    rx = 0;
    #5208
    #5208
    rx = 1;


 
end
always begin
    #1 clk = 0;
    #1 clk = 1;
end

uart uart_u(
    .clk(clk),
    .rst_p(rst),
    .uart_rx(rx),
    .uart_done(flag),
    .buffer(data),
    .data_addr(addr)


);


endmodule

module IFU(
	input
    );
endmodule

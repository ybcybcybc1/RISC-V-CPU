//****************************
//	top module of cpu core
//****************************
`include	"D:\Grade2\RISC_V\CPU\CPU.srcs\sources_1\config.v"
module cpu_top(

    );
endmodule
